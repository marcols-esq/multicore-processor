`define INST_ADDR_W 32
`define DATA_ADDR_W 32
`define REG_ADDR_W 5
`define INST_W 32
`define DATA_W 32